`include "axi_test_base.sv"
`include "axi_test_fixied.sv"
`include "axi_test_increment.sv"
`include "axi_test_wrapping.sv"
`include "axi_test_incr_4tr.sv"
`include "axi_test_wrp_4tr.sv"
`include "axi_test_unalined_tr.sv"
`include "axi_test_slave_error.sv"
